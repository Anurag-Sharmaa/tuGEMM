`timescale 1ns / 1ps


module tuGEMM_tb();

reg clk=0;
reg rst;
reg [511:0] vector_a;
reg [511:0] vector_b;

tuGEMM_8x8 uut (
clk,
rst,
vector_a,
vector_b
    );

always #5 clk = ~clk;

initial begin
 rst = 1;
 #10
 
 rst = 0;
 
// // positive values
//vector_a = 512'b00010000000011110000111000001101000011000000101100001010000010010000100000000111000001100000010100000100000000110000001000000001000100000000111100001110000011010000110000001011000010100000100100001000000001110000011000000101000001000000001100000010000000010001000000001111000011100000110100001100000010110000101000001001000010000000011100000110000001010000010000000011000000100000000100010000000011110000111000001101000011000000101100001010000010010000100000000111000001100000010100000100000000110000001000000001;

//vector_b = 512'b00000001000000100000010000000010000000100000001100000100000001010000010100000100000000110000001000000011000001000000001000000001000000010000001000000100000000100000001000000011000001000000010100000101000001000000001100000010000000110000010000000010000000010000000100000010000001000000001000000010000000110000010000000101000001010000010000000011000000100000001100000100000000100000000100000001000000100000010000000010000000100000001100000100000001010000010100000100000000110000001000000011000001000000001000000001;

// negative values
//  vector_a = 128'b00010000111100011111001000001101111101000000101111110110000010010000100011111001111110100000010100000100111111010000001011111111;
//  vector_b = 128'b11111111111111100000010011111110000000101111110111111100000001011111101100000100111111010000001011111101000001001111111000000001;

//Approx ZLCADCT
// Cameraman_txt
//vector_a = 512'b00000000000000001111111100000000000000000000000100000000000000000000000011111111000000010000000000000000000000011111111100000000000000000000000000000000111111110000000100000000000000000000000000000001111111111111111100000001000000011111111111111111000000011111111100000000000000000000000000000000000000000000000000000001000000010000000000000000111111111111111100000000000000000000000100000000111111110000000000000000000000000000000000000001000000000000000100000001000000010000000100000001000000010000000100000001;
//vector_b = 512'b11010100110101011101010111010011110100111101001111010110110101011101001111010001110100011101001011010110110101101101011011010011110101111101001111010100110100101101010111010101110101011101010111010010110101011101001011010101110101001101010011010111110101011101000011010100110100011101010111010101110101001101010111010011110101011100111111010101110101011101100111010011110110001101010111010011110100111101010011010101110101111101001011010101110101001101010111010101110100111101001111010101110101011101010011010010;


//cameraman_error
vector_a = 512'b00000000000000001111111100000000000000000000000100000000000000000000000011111111000000010000000000000000000000011111111100000000000000000000000000000000111111110000000100000000000000000000000000000001111111111111111100000001000000011111111111111111000000011111111100000000000000000000000000000000000000000000000000000001000000010000000000000000111111111111111100000000000000000000000100000000111111110000000000000000000000000000000000000001000000000000000100000001000000010000000100000001000000010000000100000001;

  vector_b = 512'b00000110000000110000011000000000111111101111111100000001000000100000001011111100111111111111110000000001000000100000000100000000000001111111111100000011111111010000000000000001000000000000001000000011000000100000001000000001111111110000000000000010000000101111101111111111111111000000000001010100010100110101010001010010111111001111011011111100111111000101100001010010010101110101010011111100111111001111110111111110010101100101000101010100010100110000000000000000111111101111111001010100010101000101001101010001;
 
 
end


endmodule
